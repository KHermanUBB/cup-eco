magic
tech sky130A
magscale 1 2
timestamp 1636601814
<< obsli1 >>
rect 1104 1377 499439 497777
<< obsm1 >>
rect 474 1368 499454 497808
<< metal2 >>
rect 2134 499200 2190 500000
rect 6458 499200 6514 500000
rect 10782 499200 10838 500000
rect 15106 499200 15162 500000
rect 19522 499200 19578 500000
rect 23846 499200 23902 500000
rect 28170 499200 28226 500000
rect 32494 499200 32550 500000
rect 36910 499200 36966 500000
rect 41234 499200 41290 500000
rect 45558 499200 45614 500000
rect 49882 499200 49938 500000
rect 54298 499200 54354 500000
rect 58622 499200 58678 500000
rect 62946 499200 63002 500000
rect 67270 499200 67326 500000
rect 71686 499200 71742 500000
rect 76010 499200 76066 500000
rect 80334 499200 80390 500000
rect 84658 499200 84714 500000
rect 89074 499200 89130 500000
rect 93398 499200 93454 500000
rect 97722 499200 97778 500000
rect 102138 499200 102194 500000
rect 106462 499200 106518 500000
rect 110786 499200 110842 500000
rect 115110 499200 115166 500000
rect 119526 499200 119582 500000
rect 123850 499200 123906 500000
rect 128174 499200 128230 500000
rect 132498 499200 132554 500000
rect 136914 499200 136970 500000
rect 141238 499200 141294 500000
rect 145562 499200 145618 500000
rect 149886 499200 149942 500000
rect 154302 499200 154358 500000
rect 158626 499200 158682 500000
rect 162950 499200 163006 500000
rect 167274 499200 167330 500000
rect 171690 499200 171746 500000
rect 176014 499200 176070 500000
rect 180338 499200 180394 500000
rect 184662 499200 184718 500000
rect 189078 499200 189134 500000
rect 193402 499200 193458 500000
rect 197726 499200 197782 500000
rect 202142 499200 202198 500000
rect 206466 499200 206522 500000
rect 210790 499200 210846 500000
rect 215114 499200 215170 500000
rect 219530 499200 219586 500000
rect 223854 499200 223910 500000
rect 228178 499200 228234 500000
rect 232502 499200 232558 500000
rect 236918 499200 236974 500000
rect 241242 499200 241298 500000
rect 245566 499200 245622 500000
rect 249890 499200 249946 500000
rect 254306 499200 254362 500000
rect 258630 499200 258686 500000
rect 262954 499200 263010 500000
rect 267278 499200 267334 500000
rect 271694 499200 271750 500000
rect 276018 499200 276074 500000
rect 280342 499200 280398 500000
rect 284666 499200 284722 500000
rect 289082 499200 289138 500000
rect 293406 499200 293462 500000
rect 297730 499200 297786 500000
rect 302146 499200 302202 500000
rect 306470 499200 306526 500000
rect 310794 499200 310850 500000
rect 315118 499200 315174 500000
rect 319534 499200 319590 500000
rect 323858 499200 323914 500000
rect 328182 499200 328238 500000
rect 332506 499200 332562 500000
rect 336922 499200 336978 500000
rect 341246 499200 341302 500000
rect 345570 499200 345626 500000
rect 349894 499200 349950 500000
rect 354310 499200 354366 500000
rect 358634 499200 358690 500000
rect 362958 499200 363014 500000
rect 367282 499200 367338 500000
rect 371698 499200 371754 500000
rect 376022 499200 376078 500000
rect 380346 499200 380402 500000
rect 384670 499200 384726 500000
rect 389086 499200 389142 500000
rect 393410 499200 393466 500000
rect 397734 499200 397790 500000
rect 402150 499200 402206 500000
rect 406474 499200 406530 500000
rect 410798 499200 410854 500000
rect 415122 499200 415178 500000
rect 419538 499200 419594 500000
rect 423862 499200 423918 500000
rect 428186 499200 428242 500000
rect 432510 499200 432566 500000
rect 436926 499200 436982 500000
rect 441250 499200 441306 500000
rect 445574 499200 445630 500000
rect 449898 499200 449954 500000
rect 454314 499200 454370 500000
rect 458638 499200 458694 500000
rect 462962 499200 463018 500000
rect 467286 499200 467342 500000
rect 471702 499200 471758 500000
rect 476026 499200 476082 500000
rect 480350 499200 480406 500000
rect 484674 499200 484730 500000
rect 489090 499200 489146 500000
rect 493414 499200 493470 500000
rect 497738 499200 497794 500000
rect 478 0 534 800
rect 1490 0 1546 800
rect 2502 0 2558 800
rect 3514 0 3570 800
rect 4526 0 4582 800
rect 5538 0 5594 800
rect 6550 0 6606 800
rect 7562 0 7618 800
rect 8574 0 8630 800
rect 9586 0 9642 800
rect 10598 0 10654 800
rect 11610 0 11666 800
rect 12622 0 12678 800
rect 13634 0 13690 800
rect 14646 0 14702 800
rect 15658 0 15714 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18694 0 18750 800
rect 19706 0 19762 800
rect 20718 0 20774 800
rect 21730 0 21786 800
rect 22742 0 22798 800
rect 23754 0 23810 800
rect 24766 0 24822 800
rect 25778 0 25834 800
rect 26790 0 26846 800
rect 27802 0 27858 800
rect 28814 0 28870 800
rect 29826 0 29882 800
rect 30838 0 30894 800
rect 31850 0 31906 800
rect 32862 0 32918 800
rect 33874 0 33930 800
rect 34886 0 34942 800
rect 35898 0 35954 800
rect 36910 0 36966 800
rect 37922 0 37978 800
rect 38934 0 38990 800
rect 39946 0 40002 800
rect 40958 0 41014 800
rect 41970 0 42026 800
rect 43074 0 43130 800
rect 44086 0 44142 800
rect 45098 0 45154 800
rect 46110 0 46166 800
rect 47122 0 47178 800
rect 48134 0 48190 800
rect 49146 0 49202 800
rect 50158 0 50214 800
rect 51170 0 51226 800
rect 52182 0 52238 800
rect 53194 0 53250 800
rect 54206 0 54262 800
rect 55218 0 55274 800
rect 56230 0 56286 800
rect 57242 0 57298 800
rect 58254 0 58310 800
rect 59266 0 59322 800
rect 60278 0 60334 800
rect 61290 0 61346 800
rect 62302 0 62358 800
rect 63314 0 63370 800
rect 64326 0 64382 800
rect 65338 0 65394 800
rect 66350 0 66406 800
rect 67362 0 67418 800
rect 68374 0 68430 800
rect 69386 0 69442 800
rect 70398 0 70454 800
rect 71410 0 71466 800
rect 72422 0 72478 800
rect 73434 0 73490 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76470 0 76526 800
rect 77482 0 77538 800
rect 78494 0 78550 800
rect 79506 0 79562 800
rect 80518 0 80574 800
rect 81530 0 81586 800
rect 82542 0 82598 800
rect 83554 0 83610 800
rect 84658 0 84714 800
rect 85670 0 85726 800
rect 86682 0 86738 800
rect 87694 0 87750 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90730 0 90786 800
rect 91742 0 91798 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94778 0 94834 800
rect 95790 0 95846 800
rect 96802 0 96858 800
rect 97814 0 97870 800
rect 98826 0 98882 800
rect 99838 0 99894 800
rect 100850 0 100906 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103886 0 103942 800
rect 104898 0 104954 800
rect 105910 0 105966 800
rect 106922 0 106978 800
rect 107934 0 107990 800
rect 108946 0 109002 800
rect 109958 0 110014 800
rect 110970 0 111026 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 114006 0 114062 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 117042 0 117098 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 121090 0 121146 800
rect 122102 0 122158 800
rect 123114 0 123170 800
rect 124126 0 124182 800
rect 125138 0 125194 800
rect 126242 0 126298 800
rect 127254 0 127310 800
rect 128266 0 128322 800
rect 129278 0 129334 800
rect 130290 0 130346 800
rect 131302 0 131358 800
rect 132314 0 132370 800
rect 133326 0 133382 800
rect 134338 0 134394 800
rect 135350 0 135406 800
rect 136362 0 136418 800
rect 137374 0 137430 800
rect 138386 0 138442 800
rect 139398 0 139454 800
rect 140410 0 140466 800
rect 141422 0 141478 800
rect 142434 0 142490 800
rect 143446 0 143502 800
rect 144458 0 144514 800
rect 145470 0 145526 800
rect 146482 0 146538 800
rect 147494 0 147550 800
rect 148506 0 148562 800
rect 149518 0 149574 800
rect 150530 0 150586 800
rect 151542 0 151598 800
rect 152554 0 152610 800
rect 153566 0 153622 800
rect 154578 0 154634 800
rect 155590 0 155646 800
rect 156602 0 156658 800
rect 157614 0 157670 800
rect 158626 0 158682 800
rect 159638 0 159694 800
rect 160650 0 160706 800
rect 161662 0 161718 800
rect 162674 0 162730 800
rect 163686 0 163742 800
rect 164698 0 164754 800
rect 165710 0 165766 800
rect 166722 0 166778 800
rect 167826 0 167882 800
rect 168838 0 168894 800
rect 169850 0 169906 800
rect 170862 0 170918 800
rect 171874 0 171930 800
rect 172886 0 172942 800
rect 173898 0 173954 800
rect 174910 0 174966 800
rect 175922 0 175978 800
rect 176934 0 176990 800
rect 177946 0 178002 800
rect 178958 0 179014 800
rect 179970 0 180026 800
rect 180982 0 181038 800
rect 181994 0 182050 800
rect 183006 0 183062 800
rect 184018 0 184074 800
rect 185030 0 185086 800
rect 186042 0 186098 800
rect 187054 0 187110 800
rect 188066 0 188122 800
rect 189078 0 189134 800
rect 190090 0 190146 800
rect 191102 0 191158 800
rect 192114 0 192170 800
rect 193126 0 193182 800
rect 194138 0 194194 800
rect 195150 0 195206 800
rect 196162 0 196218 800
rect 197174 0 197230 800
rect 198186 0 198242 800
rect 199198 0 199254 800
rect 200210 0 200266 800
rect 201222 0 201278 800
rect 202234 0 202290 800
rect 203246 0 203302 800
rect 204258 0 204314 800
rect 205270 0 205326 800
rect 206282 0 206338 800
rect 207294 0 207350 800
rect 208306 0 208362 800
rect 209410 0 209466 800
rect 210422 0 210478 800
rect 211434 0 211490 800
rect 212446 0 212502 800
rect 213458 0 213514 800
rect 214470 0 214526 800
rect 215482 0 215538 800
rect 216494 0 216550 800
rect 217506 0 217562 800
rect 218518 0 218574 800
rect 219530 0 219586 800
rect 220542 0 220598 800
rect 221554 0 221610 800
rect 222566 0 222622 800
rect 223578 0 223634 800
rect 224590 0 224646 800
rect 225602 0 225658 800
rect 226614 0 226670 800
rect 227626 0 227682 800
rect 228638 0 228694 800
rect 229650 0 229706 800
rect 230662 0 230718 800
rect 231674 0 231730 800
rect 232686 0 232742 800
rect 233698 0 233754 800
rect 234710 0 234766 800
rect 235722 0 235778 800
rect 236734 0 236790 800
rect 237746 0 237802 800
rect 238758 0 238814 800
rect 239770 0 239826 800
rect 240782 0 240838 800
rect 241794 0 241850 800
rect 242806 0 242862 800
rect 243818 0 243874 800
rect 244830 0 244886 800
rect 245842 0 245898 800
rect 246854 0 246910 800
rect 247866 0 247922 800
rect 248878 0 248934 800
rect 249890 0 249946 800
rect 250994 0 251050 800
rect 252006 0 252062 800
rect 253018 0 253074 800
rect 254030 0 254086 800
rect 255042 0 255098 800
rect 256054 0 256110 800
rect 257066 0 257122 800
rect 258078 0 258134 800
rect 259090 0 259146 800
rect 260102 0 260158 800
rect 261114 0 261170 800
rect 262126 0 262182 800
rect 263138 0 263194 800
rect 264150 0 264206 800
rect 265162 0 265218 800
rect 266174 0 266230 800
rect 267186 0 267242 800
rect 268198 0 268254 800
rect 269210 0 269266 800
rect 270222 0 270278 800
rect 271234 0 271290 800
rect 272246 0 272302 800
rect 273258 0 273314 800
rect 274270 0 274326 800
rect 275282 0 275338 800
rect 276294 0 276350 800
rect 277306 0 277362 800
rect 278318 0 278374 800
rect 279330 0 279386 800
rect 280342 0 280398 800
rect 281354 0 281410 800
rect 282366 0 282422 800
rect 283378 0 283434 800
rect 284390 0 284446 800
rect 285402 0 285458 800
rect 286414 0 286470 800
rect 287426 0 287482 800
rect 288438 0 288494 800
rect 289450 0 289506 800
rect 290462 0 290518 800
rect 291474 0 291530 800
rect 292578 0 292634 800
rect 293590 0 293646 800
rect 294602 0 294658 800
rect 295614 0 295670 800
rect 296626 0 296682 800
rect 297638 0 297694 800
rect 298650 0 298706 800
rect 299662 0 299718 800
rect 300674 0 300730 800
rect 301686 0 301742 800
rect 302698 0 302754 800
rect 303710 0 303766 800
rect 304722 0 304778 800
rect 305734 0 305790 800
rect 306746 0 306802 800
rect 307758 0 307814 800
rect 308770 0 308826 800
rect 309782 0 309838 800
rect 310794 0 310850 800
rect 311806 0 311862 800
rect 312818 0 312874 800
rect 313830 0 313886 800
rect 314842 0 314898 800
rect 315854 0 315910 800
rect 316866 0 316922 800
rect 317878 0 317934 800
rect 318890 0 318946 800
rect 319902 0 319958 800
rect 320914 0 320970 800
rect 321926 0 321982 800
rect 322938 0 322994 800
rect 323950 0 324006 800
rect 324962 0 325018 800
rect 325974 0 326030 800
rect 326986 0 327042 800
rect 327998 0 328054 800
rect 329010 0 329066 800
rect 330022 0 330078 800
rect 331034 0 331090 800
rect 332046 0 332102 800
rect 333058 0 333114 800
rect 334162 0 334218 800
rect 335174 0 335230 800
rect 336186 0 336242 800
rect 337198 0 337254 800
rect 338210 0 338266 800
rect 339222 0 339278 800
rect 340234 0 340290 800
rect 341246 0 341302 800
rect 342258 0 342314 800
rect 343270 0 343326 800
rect 344282 0 344338 800
rect 345294 0 345350 800
rect 346306 0 346362 800
rect 347318 0 347374 800
rect 348330 0 348386 800
rect 349342 0 349398 800
rect 350354 0 350410 800
rect 351366 0 351422 800
rect 352378 0 352434 800
rect 353390 0 353446 800
rect 354402 0 354458 800
rect 355414 0 355470 800
rect 356426 0 356482 800
rect 357438 0 357494 800
rect 358450 0 358506 800
rect 359462 0 359518 800
rect 360474 0 360530 800
rect 361486 0 361542 800
rect 362498 0 362554 800
rect 363510 0 363566 800
rect 364522 0 364578 800
rect 365534 0 365590 800
rect 366546 0 366602 800
rect 367558 0 367614 800
rect 368570 0 368626 800
rect 369582 0 369638 800
rect 370594 0 370650 800
rect 371606 0 371662 800
rect 372618 0 372674 800
rect 373630 0 373686 800
rect 374642 0 374698 800
rect 375746 0 375802 800
rect 376758 0 376814 800
rect 377770 0 377826 800
rect 378782 0 378838 800
rect 379794 0 379850 800
rect 380806 0 380862 800
rect 381818 0 381874 800
rect 382830 0 382886 800
rect 383842 0 383898 800
rect 384854 0 384910 800
rect 385866 0 385922 800
rect 386878 0 386934 800
rect 387890 0 387946 800
rect 388902 0 388958 800
rect 389914 0 389970 800
rect 390926 0 390982 800
rect 391938 0 391994 800
rect 392950 0 393006 800
rect 393962 0 394018 800
rect 394974 0 395030 800
rect 395986 0 396042 800
rect 396998 0 397054 800
rect 398010 0 398066 800
rect 399022 0 399078 800
rect 400034 0 400090 800
rect 401046 0 401102 800
rect 402058 0 402114 800
rect 403070 0 403126 800
rect 404082 0 404138 800
rect 405094 0 405150 800
rect 406106 0 406162 800
rect 407118 0 407174 800
rect 408130 0 408186 800
rect 409142 0 409198 800
rect 410154 0 410210 800
rect 411166 0 411222 800
rect 412178 0 412234 800
rect 413190 0 413246 800
rect 414202 0 414258 800
rect 415214 0 415270 800
rect 416226 0 416282 800
rect 417330 0 417386 800
rect 418342 0 418398 800
rect 419354 0 419410 800
rect 420366 0 420422 800
rect 421378 0 421434 800
rect 422390 0 422446 800
rect 423402 0 423458 800
rect 424414 0 424470 800
rect 425426 0 425482 800
rect 426438 0 426494 800
rect 427450 0 427506 800
rect 428462 0 428518 800
rect 429474 0 429530 800
rect 430486 0 430542 800
rect 431498 0 431554 800
rect 432510 0 432566 800
rect 433522 0 433578 800
rect 434534 0 434590 800
rect 435546 0 435602 800
rect 436558 0 436614 800
rect 437570 0 437626 800
rect 438582 0 438638 800
rect 439594 0 439650 800
rect 440606 0 440662 800
rect 441618 0 441674 800
rect 442630 0 442686 800
rect 443642 0 443698 800
rect 444654 0 444710 800
rect 445666 0 445722 800
rect 446678 0 446734 800
rect 447690 0 447746 800
rect 448702 0 448758 800
rect 449714 0 449770 800
rect 450726 0 450782 800
rect 451738 0 451794 800
rect 452750 0 452806 800
rect 453762 0 453818 800
rect 454774 0 454830 800
rect 455786 0 455842 800
rect 456798 0 456854 800
rect 457810 0 457866 800
rect 458914 0 458970 800
rect 459926 0 459982 800
rect 460938 0 460994 800
rect 461950 0 462006 800
rect 462962 0 463018 800
rect 463974 0 464030 800
rect 464986 0 465042 800
rect 465998 0 466054 800
rect 467010 0 467066 800
rect 468022 0 468078 800
rect 469034 0 469090 800
rect 470046 0 470102 800
rect 471058 0 471114 800
rect 472070 0 472126 800
rect 473082 0 473138 800
rect 474094 0 474150 800
rect 475106 0 475162 800
rect 476118 0 476174 800
rect 477130 0 477186 800
rect 478142 0 478198 800
rect 479154 0 479210 800
rect 480166 0 480222 800
rect 481178 0 481234 800
rect 482190 0 482246 800
rect 483202 0 483258 800
rect 484214 0 484270 800
rect 485226 0 485282 800
rect 486238 0 486294 800
rect 487250 0 487306 800
rect 488262 0 488318 800
rect 489274 0 489330 800
rect 490286 0 490342 800
rect 491298 0 491354 800
rect 492310 0 492366 800
rect 493322 0 493378 800
rect 494334 0 494390 800
rect 495346 0 495402 800
rect 496358 0 496414 800
rect 497370 0 497426 800
rect 498382 0 498438 800
rect 499394 0 499450 800
<< obsm2 >>
rect 480 499144 2078 499338
rect 2246 499144 6402 499338
rect 6570 499144 10726 499338
rect 10894 499144 15050 499338
rect 15218 499144 19466 499338
rect 19634 499144 23790 499338
rect 23958 499144 28114 499338
rect 28282 499144 32438 499338
rect 32606 499144 36854 499338
rect 37022 499144 41178 499338
rect 41346 499144 45502 499338
rect 45670 499144 49826 499338
rect 49994 499144 54242 499338
rect 54410 499144 58566 499338
rect 58734 499144 62890 499338
rect 63058 499144 67214 499338
rect 67382 499144 71630 499338
rect 71798 499144 75954 499338
rect 76122 499144 80278 499338
rect 80446 499144 84602 499338
rect 84770 499144 89018 499338
rect 89186 499144 93342 499338
rect 93510 499144 97666 499338
rect 97834 499144 102082 499338
rect 102250 499144 106406 499338
rect 106574 499144 110730 499338
rect 110898 499144 115054 499338
rect 115222 499144 119470 499338
rect 119638 499144 123794 499338
rect 123962 499144 128118 499338
rect 128286 499144 132442 499338
rect 132610 499144 136858 499338
rect 137026 499144 141182 499338
rect 141350 499144 145506 499338
rect 145674 499144 149830 499338
rect 149998 499144 154246 499338
rect 154414 499144 158570 499338
rect 158738 499144 162894 499338
rect 163062 499144 167218 499338
rect 167386 499144 171634 499338
rect 171802 499144 175958 499338
rect 176126 499144 180282 499338
rect 180450 499144 184606 499338
rect 184774 499144 189022 499338
rect 189190 499144 193346 499338
rect 193514 499144 197670 499338
rect 197838 499144 202086 499338
rect 202254 499144 206410 499338
rect 206578 499144 210734 499338
rect 210902 499144 215058 499338
rect 215226 499144 219474 499338
rect 219642 499144 223798 499338
rect 223966 499144 228122 499338
rect 228290 499144 232446 499338
rect 232614 499144 236862 499338
rect 237030 499144 241186 499338
rect 241354 499144 245510 499338
rect 245678 499144 249834 499338
rect 250002 499144 254250 499338
rect 254418 499144 258574 499338
rect 258742 499144 262898 499338
rect 263066 499144 267222 499338
rect 267390 499144 271638 499338
rect 271806 499144 275962 499338
rect 276130 499144 280286 499338
rect 280454 499144 284610 499338
rect 284778 499144 289026 499338
rect 289194 499144 293350 499338
rect 293518 499144 297674 499338
rect 297842 499144 302090 499338
rect 302258 499144 306414 499338
rect 306582 499144 310738 499338
rect 310906 499144 315062 499338
rect 315230 499144 319478 499338
rect 319646 499144 323802 499338
rect 323970 499144 328126 499338
rect 328294 499144 332450 499338
rect 332618 499144 336866 499338
rect 337034 499144 341190 499338
rect 341358 499144 345514 499338
rect 345682 499144 349838 499338
rect 350006 499144 354254 499338
rect 354422 499144 358578 499338
rect 358746 499144 362902 499338
rect 363070 499144 367226 499338
rect 367394 499144 371642 499338
rect 371810 499144 375966 499338
rect 376134 499144 380290 499338
rect 380458 499144 384614 499338
rect 384782 499144 389030 499338
rect 389198 499144 393354 499338
rect 393522 499144 397678 499338
rect 397846 499144 402094 499338
rect 402262 499144 406418 499338
rect 406586 499144 410742 499338
rect 410910 499144 415066 499338
rect 415234 499144 419482 499338
rect 419650 499144 423806 499338
rect 423974 499144 428130 499338
rect 428298 499144 432454 499338
rect 432622 499144 436870 499338
rect 437038 499144 441194 499338
rect 441362 499144 445518 499338
rect 445686 499144 449842 499338
rect 450010 499144 454258 499338
rect 454426 499144 458582 499338
rect 458750 499144 462906 499338
rect 463074 499144 467230 499338
rect 467398 499144 471646 499338
rect 471814 499144 475970 499338
rect 476138 499144 480294 499338
rect 480462 499144 484618 499338
rect 484786 499144 489034 499338
rect 489202 499144 493358 499338
rect 493526 499144 497682 499338
rect 497850 499144 499448 499338
rect 480 856 499448 499144
rect 590 734 1434 856
rect 1602 734 2446 856
rect 2614 734 3458 856
rect 3626 734 4470 856
rect 4638 734 5482 856
rect 5650 734 6494 856
rect 6662 734 7506 856
rect 7674 734 8518 856
rect 8686 734 9530 856
rect 9698 734 10542 856
rect 10710 734 11554 856
rect 11722 734 12566 856
rect 12734 734 13578 856
rect 13746 734 14590 856
rect 14758 734 15602 856
rect 15770 734 16614 856
rect 16782 734 17626 856
rect 17794 734 18638 856
rect 18806 734 19650 856
rect 19818 734 20662 856
rect 20830 734 21674 856
rect 21842 734 22686 856
rect 22854 734 23698 856
rect 23866 734 24710 856
rect 24878 734 25722 856
rect 25890 734 26734 856
rect 26902 734 27746 856
rect 27914 734 28758 856
rect 28926 734 29770 856
rect 29938 734 30782 856
rect 30950 734 31794 856
rect 31962 734 32806 856
rect 32974 734 33818 856
rect 33986 734 34830 856
rect 34998 734 35842 856
rect 36010 734 36854 856
rect 37022 734 37866 856
rect 38034 734 38878 856
rect 39046 734 39890 856
rect 40058 734 40902 856
rect 41070 734 41914 856
rect 42082 734 43018 856
rect 43186 734 44030 856
rect 44198 734 45042 856
rect 45210 734 46054 856
rect 46222 734 47066 856
rect 47234 734 48078 856
rect 48246 734 49090 856
rect 49258 734 50102 856
rect 50270 734 51114 856
rect 51282 734 52126 856
rect 52294 734 53138 856
rect 53306 734 54150 856
rect 54318 734 55162 856
rect 55330 734 56174 856
rect 56342 734 57186 856
rect 57354 734 58198 856
rect 58366 734 59210 856
rect 59378 734 60222 856
rect 60390 734 61234 856
rect 61402 734 62246 856
rect 62414 734 63258 856
rect 63426 734 64270 856
rect 64438 734 65282 856
rect 65450 734 66294 856
rect 66462 734 67306 856
rect 67474 734 68318 856
rect 68486 734 69330 856
rect 69498 734 70342 856
rect 70510 734 71354 856
rect 71522 734 72366 856
rect 72534 734 73378 856
rect 73546 734 74390 856
rect 74558 734 75402 856
rect 75570 734 76414 856
rect 76582 734 77426 856
rect 77594 734 78438 856
rect 78606 734 79450 856
rect 79618 734 80462 856
rect 80630 734 81474 856
rect 81642 734 82486 856
rect 82654 734 83498 856
rect 83666 734 84602 856
rect 84770 734 85614 856
rect 85782 734 86626 856
rect 86794 734 87638 856
rect 87806 734 88650 856
rect 88818 734 89662 856
rect 89830 734 90674 856
rect 90842 734 91686 856
rect 91854 734 92698 856
rect 92866 734 93710 856
rect 93878 734 94722 856
rect 94890 734 95734 856
rect 95902 734 96746 856
rect 96914 734 97758 856
rect 97926 734 98770 856
rect 98938 734 99782 856
rect 99950 734 100794 856
rect 100962 734 101806 856
rect 101974 734 102818 856
rect 102986 734 103830 856
rect 103998 734 104842 856
rect 105010 734 105854 856
rect 106022 734 106866 856
rect 107034 734 107878 856
rect 108046 734 108890 856
rect 109058 734 109902 856
rect 110070 734 110914 856
rect 111082 734 111926 856
rect 112094 734 112938 856
rect 113106 734 113950 856
rect 114118 734 114962 856
rect 115130 734 115974 856
rect 116142 734 116986 856
rect 117154 734 117998 856
rect 118166 734 119010 856
rect 119178 734 120022 856
rect 120190 734 121034 856
rect 121202 734 122046 856
rect 122214 734 123058 856
rect 123226 734 124070 856
rect 124238 734 125082 856
rect 125250 734 126186 856
rect 126354 734 127198 856
rect 127366 734 128210 856
rect 128378 734 129222 856
rect 129390 734 130234 856
rect 130402 734 131246 856
rect 131414 734 132258 856
rect 132426 734 133270 856
rect 133438 734 134282 856
rect 134450 734 135294 856
rect 135462 734 136306 856
rect 136474 734 137318 856
rect 137486 734 138330 856
rect 138498 734 139342 856
rect 139510 734 140354 856
rect 140522 734 141366 856
rect 141534 734 142378 856
rect 142546 734 143390 856
rect 143558 734 144402 856
rect 144570 734 145414 856
rect 145582 734 146426 856
rect 146594 734 147438 856
rect 147606 734 148450 856
rect 148618 734 149462 856
rect 149630 734 150474 856
rect 150642 734 151486 856
rect 151654 734 152498 856
rect 152666 734 153510 856
rect 153678 734 154522 856
rect 154690 734 155534 856
rect 155702 734 156546 856
rect 156714 734 157558 856
rect 157726 734 158570 856
rect 158738 734 159582 856
rect 159750 734 160594 856
rect 160762 734 161606 856
rect 161774 734 162618 856
rect 162786 734 163630 856
rect 163798 734 164642 856
rect 164810 734 165654 856
rect 165822 734 166666 856
rect 166834 734 167770 856
rect 167938 734 168782 856
rect 168950 734 169794 856
rect 169962 734 170806 856
rect 170974 734 171818 856
rect 171986 734 172830 856
rect 172998 734 173842 856
rect 174010 734 174854 856
rect 175022 734 175866 856
rect 176034 734 176878 856
rect 177046 734 177890 856
rect 178058 734 178902 856
rect 179070 734 179914 856
rect 180082 734 180926 856
rect 181094 734 181938 856
rect 182106 734 182950 856
rect 183118 734 183962 856
rect 184130 734 184974 856
rect 185142 734 185986 856
rect 186154 734 186998 856
rect 187166 734 188010 856
rect 188178 734 189022 856
rect 189190 734 190034 856
rect 190202 734 191046 856
rect 191214 734 192058 856
rect 192226 734 193070 856
rect 193238 734 194082 856
rect 194250 734 195094 856
rect 195262 734 196106 856
rect 196274 734 197118 856
rect 197286 734 198130 856
rect 198298 734 199142 856
rect 199310 734 200154 856
rect 200322 734 201166 856
rect 201334 734 202178 856
rect 202346 734 203190 856
rect 203358 734 204202 856
rect 204370 734 205214 856
rect 205382 734 206226 856
rect 206394 734 207238 856
rect 207406 734 208250 856
rect 208418 734 209354 856
rect 209522 734 210366 856
rect 210534 734 211378 856
rect 211546 734 212390 856
rect 212558 734 213402 856
rect 213570 734 214414 856
rect 214582 734 215426 856
rect 215594 734 216438 856
rect 216606 734 217450 856
rect 217618 734 218462 856
rect 218630 734 219474 856
rect 219642 734 220486 856
rect 220654 734 221498 856
rect 221666 734 222510 856
rect 222678 734 223522 856
rect 223690 734 224534 856
rect 224702 734 225546 856
rect 225714 734 226558 856
rect 226726 734 227570 856
rect 227738 734 228582 856
rect 228750 734 229594 856
rect 229762 734 230606 856
rect 230774 734 231618 856
rect 231786 734 232630 856
rect 232798 734 233642 856
rect 233810 734 234654 856
rect 234822 734 235666 856
rect 235834 734 236678 856
rect 236846 734 237690 856
rect 237858 734 238702 856
rect 238870 734 239714 856
rect 239882 734 240726 856
rect 240894 734 241738 856
rect 241906 734 242750 856
rect 242918 734 243762 856
rect 243930 734 244774 856
rect 244942 734 245786 856
rect 245954 734 246798 856
rect 246966 734 247810 856
rect 247978 734 248822 856
rect 248990 734 249834 856
rect 250002 734 250938 856
rect 251106 734 251950 856
rect 252118 734 252962 856
rect 253130 734 253974 856
rect 254142 734 254986 856
rect 255154 734 255998 856
rect 256166 734 257010 856
rect 257178 734 258022 856
rect 258190 734 259034 856
rect 259202 734 260046 856
rect 260214 734 261058 856
rect 261226 734 262070 856
rect 262238 734 263082 856
rect 263250 734 264094 856
rect 264262 734 265106 856
rect 265274 734 266118 856
rect 266286 734 267130 856
rect 267298 734 268142 856
rect 268310 734 269154 856
rect 269322 734 270166 856
rect 270334 734 271178 856
rect 271346 734 272190 856
rect 272358 734 273202 856
rect 273370 734 274214 856
rect 274382 734 275226 856
rect 275394 734 276238 856
rect 276406 734 277250 856
rect 277418 734 278262 856
rect 278430 734 279274 856
rect 279442 734 280286 856
rect 280454 734 281298 856
rect 281466 734 282310 856
rect 282478 734 283322 856
rect 283490 734 284334 856
rect 284502 734 285346 856
rect 285514 734 286358 856
rect 286526 734 287370 856
rect 287538 734 288382 856
rect 288550 734 289394 856
rect 289562 734 290406 856
rect 290574 734 291418 856
rect 291586 734 292522 856
rect 292690 734 293534 856
rect 293702 734 294546 856
rect 294714 734 295558 856
rect 295726 734 296570 856
rect 296738 734 297582 856
rect 297750 734 298594 856
rect 298762 734 299606 856
rect 299774 734 300618 856
rect 300786 734 301630 856
rect 301798 734 302642 856
rect 302810 734 303654 856
rect 303822 734 304666 856
rect 304834 734 305678 856
rect 305846 734 306690 856
rect 306858 734 307702 856
rect 307870 734 308714 856
rect 308882 734 309726 856
rect 309894 734 310738 856
rect 310906 734 311750 856
rect 311918 734 312762 856
rect 312930 734 313774 856
rect 313942 734 314786 856
rect 314954 734 315798 856
rect 315966 734 316810 856
rect 316978 734 317822 856
rect 317990 734 318834 856
rect 319002 734 319846 856
rect 320014 734 320858 856
rect 321026 734 321870 856
rect 322038 734 322882 856
rect 323050 734 323894 856
rect 324062 734 324906 856
rect 325074 734 325918 856
rect 326086 734 326930 856
rect 327098 734 327942 856
rect 328110 734 328954 856
rect 329122 734 329966 856
rect 330134 734 330978 856
rect 331146 734 331990 856
rect 332158 734 333002 856
rect 333170 734 334106 856
rect 334274 734 335118 856
rect 335286 734 336130 856
rect 336298 734 337142 856
rect 337310 734 338154 856
rect 338322 734 339166 856
rect 339334 734 340178 856
rect 340346 734 341190 856
rect 341358 734 342202 856
rect 342370 734 343214 856
rect 343382 734 344226 856
rect 344394 734 345238 856
rect 345406 734 346250 856
rect 346418 734 347262 856
rect 347430 734 348274 856
rect 348442 734 349286 856
rect 349454 734 350298 856
rect 350466 734 351310 856
rect 351478 734 352322 856
rect 352490 734 353334 856
rect 353502 734 354346 856
rect 354514 734 355358 856
rect 355526 734 356370 856
rect 356538 734 357382 856
rect 357550 734 358394 856
rect 358562 734 359406 856
rect 359574 734 360418 856
rect 360586 734 361430 856
rect 361598 734 362442 856
rect 362610 734 363454 856
rect 363622 734 364466 856
rect 364634 734 365478 856
rect 365646 734 366490 856
rect 366658 734 367502 856
rect 367670 734 368514 856
rect 368682 734 369526 856
rect 369694 734 370538 856
rect 370706 734 371550 856
rect 371718 734 372562 856
rect 372730 734 373574 856
rect 373742 734 374586 856
rect 374754 734 375690 856
rect 375858 734 376702 856
rect 376870 734 377714 856
rect 377882 734 378726 856
rect 378894 734 379738 856
rect 379906 734 380750 856
rect 380918 734 381762 856
rect 381930 734 382774 856
rect 382942 734 383786 856
rect 383954 734 384798 856
rect 384966 734 385810 856
rect 385978 734 386822 856
rect 386990 734 387834 856
rect 388002 734 388846 856
rect 389014 734 389858 856
rect 390026 734 390870 856
rect 391038 734 391882 856
rect 392050 734 392894 856
rect 393062 734 393906 856
rect 394074 734 394918 856
rect 395086 734 395930 856
rect 396098 734 396942 856
rect 397110 734 397954 856
rect 398122 734 398966 856
rect 399134 734 399978 856
rect 400146 734 400990 856
rect 401158 734 402002 856
rect 402170 734 403014 856
rect 403182 734 404026 856
rect 404194 734 405038 856
rect 405206 734 406050 856
rect 406218 734 407062 856
rect 407230 734 408074 856
rect 408242 734 409086 856
rect 409254 734 410098 856
rect 410266 734 411110 856
rect 411278 734 412122 856
rect 412290 734 413134 856
rect 413302 734 414146 856
rect 414314 734 415158 856
rect 415326 734 416170 856
rect 416338 734 417274 856
rect 417442 734 418286 856
rect 418454 734 419298 856
rect 419466 734 420310 856
rect 420478 734 421322 856
rect 421490 734 422334 856
rect 422502 734 423346 856
rect 423514 734 424358 856
rect 424526 734 425370 856
rect 425538 734 426382 856
rect 426550 734 427394 856
rect 427562 734 428406 856
rect 428574 734 429418 856
rect 429586 734 430430 856
rect 430598 734 431442 856
rect 431610 734 432454 856
rect 432622 734 433466 856
rect 433634 734 434478 856
rect 434646 734 435490 856
rect 435658 734 436502 856
rect 436670 734 437514 856
rect 437682 734 438526 856
rect 438694 734 439538 856
rect 439706 734 440550 856
rect 440718 734 441562 856
rect 441730 734 442574 856
rect 442742 734 443586 856
rect 443754 734 444598 856
rect 444766 734 445610 856
rect 445778 734 446622 856
rect 446790 734 447634 856
rect 447802 734 448646 856
rect 448814 734 449658 856
rect 449826 734 450670 856
rect 450838 734 451682 856
rect 451850 734 452694 856
rect 452862 734 453706 856
rect 453874 734 454718 856
rect 454886 734 455730 856
rect 455898 734 456742 856
rect 456910 734 457754 856
rect 457922 734 458858 856
rect 459026 734 459870 856
rect 460038 734 460882 856
rect 461050 734 461894 856
rect 462062 734 462906 856
rect 463074 734 463918 856
rect 464086 734 464930 856
rect 465098 734 465942 856
rect 466110 734 466954 856
rect 467122 734 467966 856
rect 468134 734 468978 856
rect 469146 734 469990 856
rect 470158 734 471002 856
rect 471170 734 472014 856
rect 472182 734 473026 856
rect 473194 734 474038 856
rect 474206 734 475050 856
rect 475218 734 476062 856
rect 476230 734 477074 856
rect 477242 734 478086 856
rect 478254 734 479098 856
rect 479266 734 480110 856
rect 480278 734 481122 856
rect 481290 734 482134 856
rect 482302 734 483146 856
rect 483314 734 484158 856
rect 484326 734 485170 856
rect 485338 734 486182 856
rect 486350 734 487194 856
rect 487362 734 488206 856
rect 488374 734 489218 856
rect 489386 734 490230 856
rect 490398 734 491242 856
rect 491410 734 492254 856
rect 492422 734 493266 856
rect 493434 734 494278 856
rect 494446 734 495290 856
rect 495458 734 496302 856
rect 496470 734 497314 856
rect 497482 734 498326 856
rect 498494 734 499338 856
<< metal3 >>
rect 499200 249976 500000 250096
<< obsm3 >>
rect 4208 2143 496048 497793
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
rect 34928 2128 35248 497808
rect 50288 2128 50608 497808
rect 65648 2128 65968 497808
rect 81008 2128 81328 497808
rect 96368 2128 96688 497808
rect 111728 2128 112048 497808
rect 127088 2128 127408 497808
rect 142448 2128 142768 497808
rect 157808 2128 158128 497808
rect 173168 2128 173488 497808
rect 188528 2128 188848 497808
rect 203888 2128 204208 497808
rect 219248 2128 219568 497808
rect 234608 2128 234928 497808
rect 249968 2128 250288 497808
rect 265328 2128 265648 497808
rect 280688 2128 281008 497808
rect 296048 2128 296368 497808
rect 311408 2128 311728 497808
rect 326768 2128 327088 497808
rect 342128 2128 342448 497808
rect 357488 2128 357808 497808
rect 372848 2128 373168 497808
rect 388208 2128 388528 497808
rect 403568 2128 403888 497808
rect 418928 2128 419248 497808
rect 434288 2128 434608 497808
rect 449648 2128 449968 497808
rect 465008 2128 465328 497808
rect 480368 2128 480688 497808
rect 495728 2128 496048 497808
<< obsm4 >>
rect 35387 60283 50208 313309
rect 50688 60283 65568 313309
rect 66048 60283 80928 313309
rect 81408 60283 96288 313309
rect 96768 60283 111648 313309
rect 112128 60283 127008 313309
rect 127488 60283 142368 313309
rect 142848 60283 157728 313309
rect 158208 60283 173088 313309
rect 173568 60283 188448 313309
rect 188928 60283 203808 313309
rect 204288 60283 219168 313309
rect 219648 60283 234528 313309
rect 235008 60283 249888 313309
rect 250368 60283 265248 313309
rect 265728 60283 280608 313309
rect 281088 60283 295968 313309
rect 296448 60283 311328 313309
rect 311808 60283 326688 313309
rect 327168 60283 342048 313309
rect 342528 60283 357408 313309
rect 357888 60283 358373 313309
<< labels >>
rlabel metal2 s 2134 499200 2190 500000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 132498 499200 132554 500000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 145562 499200 145618 500000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 158626 499200 158682 500000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 171690 499200 171746 500000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 184662 499200 184718 500000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 197726 499200 197782 500000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 210790 499200 210846 500000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 223854 499200 223910 500000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 236918 499200 236974 500000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 249890 499200 249946 500000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 15106 499200 15162 500000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 262954 499200 263010 500000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 276018 499200 276074 500000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 289082 499200 289138 500000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 302146 499200 302202 500000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 315118 499200 315174 500000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 328182 499200 328238 500000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 341246 499200 341302 500000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 354310 499200 354366 500000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 367282 499200 367338 500000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 380346 499200 380402 500000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 28170 499200 28226 500000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 393410 499200 393466 500000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 406474 499200 406530 500000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 419538 499200 419594 500000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 432510 499200 432566 500000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 445574 499200 445630 500000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 458638 499200 458694 500000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 471702 499200 471758 500000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 484674 499200 484730 500000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 41234 499200 41290 500000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 54298 499200 54354 500000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 67270 499200 67326 500000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 80334 499200 80390 500000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 93398 499200 93454 500000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 106462 499200 106518 500000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 119526 499200 119582 500000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 499200 6514 500000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 136914 499200 136970 500000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 149886 499200 149942 500000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 162950 499200 163006 500000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 176014 499200 176070 500000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 189078 499200 189134 500000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 202142 499200 202198 500000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 215114 499200 215170 500000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 228178 499200 228234 500000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 241242 499200 241298 500000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 254306 499200 254362 500000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 19522 499200 19578 500000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 267278 499200 267334 500000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 280342 499200 280398 500000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 293406 499200 293462 500000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 306470 499200 306526 500000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 319534 499200 319590 500000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 332506 499200 332562 500000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 345570 499200 345626 500000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 358634 499200 358690 500000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 371698 499200 371754 500000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 384670 499200 384726 500000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 32494 499200 32550 500000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 397734 499200 397790 500000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 410798 499200 410854 500000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 423862 499200 423918 500000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 436926 499200 436982 500000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 449898 499200 449954 500000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 462962 499200 463018 500000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 476026 499200 476082 500000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 489090 499200 489146 500000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 45558 499200 45614 500000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 58622 499200 58678 500000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 71686 499200 71742 500000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 84658 499200 84714 500000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 97722 499200 97778 500000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 110786 499200 110842 500000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 123850 499200 123906 500000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 10782 499200 10838 500000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 141238 499200 141294 500000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 154302 499200 154358 500000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 167274 499200 167330 500000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 180338 499200 180394 500000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 193402 499200 193458 500000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 206466 499200 206522 500000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 219530 499200 219586 500000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 232502 499200 232558 500000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 245566 499200 245622 500000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 258630 499200 258686 500000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 23846 499200 23902 500000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 271694 499200 271750 500000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 284666 499200 284722 500000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 297730 499200 297786 500000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 310794 499200 310850 500000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 323858 499200 323914 500000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 336922 499200 336978 500000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 349894 499200 349950 500000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 362958 499200 363014 500000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 376022 499200 376078 500000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 389086 499200 389142 500000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 36910 499200 36966 500000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 402150 499200 402206 500000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 415122 499200 415178 500000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 428186 499200 428242 500000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 441250 499200 441306 500000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 454314 499200 454370 500000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 467286 499200 467342 500000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 480350 499200 480406 500000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 493414 499200 493470 500000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 49882 499200 49938 500000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 62946 499200 63002 500000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 76010 499200 76066 500000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 89074 499200 89130 500000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 102138 499200 102194 500000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 115110 499200 115166 500000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 128174 499200 128230 500000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 497370 0 497426 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 498382 0 498438 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 499394 0 499450 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 412178 0 412234 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 415214 0 415270 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 418342 0 418398 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 421378 0 421434 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 424414 0 424470 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 427450 0 427506 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 430486 0 430542 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 433522 0 433578 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 436558 0 436614 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 439594 0 439650 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 442630 0 442686 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 445666 0 445722 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 448702 0 448758 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 451738 0 451794 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 454774 0 454830 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 457810 0 457866 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 460938 0 460994 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 463974 0 464030 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 467010 0 467066 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 470046 0 470102 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 473082 0 473138 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 476118 0 476174 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 479154 0 479210 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 482190 0 482246 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 485226 0 485282 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 488262 0 488318 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 491298 0 491354 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 494334 0 494390 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 156602 0 156658 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 162674 0 162730 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 174910 0 174966 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 177946 0 178002 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 187054 0 187110 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 193126 0 193182 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 232686 0 232742 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 250994 0 251050 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 257066 0 257122 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 272246 0 272302 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 275282 0 275338 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 278318 0 278374 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 284390 0 284446 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 287426 0 287482 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 290462 0 290518 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 293590 0 293646 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 296626 0 296682 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 299662 0 299718 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 305734 0 305790 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 308770 0 308826 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 314842 0 314898 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 317878 0 317934 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 320914 0 320970 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 326986 0 327042 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 330022 0 330078 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 333058 0 333114 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 339222 0 339278 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 342258 0 342314 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 345294 0 345350 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 348330 0 348386 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 351366 0 351422 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 354402 0 354458 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 360474 0 360530 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 363510 0 363566 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 366546 0 366602 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 369582 0 369638 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 372618 0 372674 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 375746 0 375802 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 378782 0 378838 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 381818 0 381874 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 384854 0 384910 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 387890 0 387946 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 390926 0 390982 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 393962 0 394018 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 396998 0 397054 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 400034 0 400090 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 406106 0 406162 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 409142 0 409198 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 413190 0 413246 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 416226 0 416282 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 419354 0 419410 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 422390 0 422446 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 425426 0 425482 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 428462 0 428518 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 431498 0 431554 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 434534 0 434590 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 437570 0 437626 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 440606 0 440662 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 443642 0 443698 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 446678 0 446734 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 449714 0 449770 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 452750 0 452806 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 455786 0 455842 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 458914 0 458970 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 461950 0 462006 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 464986 0 465042 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 468022 0 468078 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 471058 0 471114 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 474094 0 474150 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 477130 0 477186 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 480166 0 480222 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 483202 0 483258 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 486238 0 486294 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 489274 0 489330 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 492310 0 492366 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 495346 0 495402 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 166722 0 166778 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 169850 0 169906 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 178958 0 179014 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 181994 0 182050 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 185030 0 185086 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 188066 0 188122 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 191102 0 191158 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 197174 0 197230 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 203246 0 203302 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 212446 0 212502 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 215482 0 215538 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 218518 0 218574 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 224590 0 224646 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 227626 0 227682 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 230662 0 230718 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 236734 0 236790 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 239770 0 239826 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 242806 0 242862 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 252006 0 252062 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 255042 0 255098 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 258078 0 258134 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 261114 0 261170 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 264150 0 264206 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 267186 0 267242 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 270222 0 270278 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 273258 0 273314 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 279330 0 279386 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 282366 0 282422 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 285402 0 285458 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 288438 0 288494 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 291474 0 291530 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 294602 0 294658 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 297638 0 297694 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 300674 0 300730 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 303710 0 303766 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 306746 0 306802 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 309782 0 309838 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 312818 0 312874 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 315854 0 315910 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 318890 0 318946 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 321926 0 321982 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 324962 0 325018 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 327998 0 328054 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 331034 0 331090 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 334162 0 334218 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 337198 0 337254 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 340234 0 340290 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 343270 0 343326 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 346306 0 346362 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 349342 0 349398 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 352378 0 352434 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 355414 0 355470 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 358450 0 358506 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 361486 0 361542 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 364522 0 364578 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 367558 0 367614 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 370594 0 370650 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 373630 0 373686 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 376758 0 376814 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 379794 0 379850 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 382830 0 382886 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 385866 0 385922 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 388902 0 388958 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 391938 0 391994 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 394974 0 395030 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 398010 0 398066 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 401046 0 401102 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 404082 0 404138 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 407118 0 407174 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 410154 0 410210 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 414202 0 414258 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 417330 0 417386 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 420366 0 420422 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 423402 0 423458 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 426438 0 426494 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 429474 0 429530 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 432510 0 432566 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 435546 0 435602 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 438582 0 438638 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 441618 0 441674 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 444654 0 444710 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 447690 0 447746 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 450726 0 450782 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 453762 0 453818 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 456798 0 456854 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 459926 0 459982 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 462962 0 463018 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 465998 0 466054 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 469034 0 469090 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 472070 0 472126 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 475106 0 475162 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 478142 0 478198 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 481178 0 481234 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 484214 0 484270 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 487250 0 487306 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 490286 0 490342 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 493322 0 493378 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 496358 0 496414 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 176934 0 176990 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 183006 0 183062 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 207294 0 207350 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 210422 0 210478 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 219530 0 219586 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 231674 0 231730 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 240782 0 240838 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 246854 0 246910 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 249890 0 249946 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 256054 0 256110 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 259090 0 259146 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 268198 0 268254 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 271234 0 271290 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 277306 0 277362 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 286414 0 286470 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 295614 0 295670 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 298650 0 298706 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 304722 0 304778 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 310794 0 310850 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 319902 0 319958 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 325974 0 326030 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 329010 0 329066 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 332046 0 332102 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 335174 0 335230 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 338210 0 338266 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 341246 0 341302 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 344282 0 344338 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 347318 0 347374 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 350354 0 350410 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 353390 0 353446 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 359462 0 359518 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 368570 0 368626 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 371606 0 371662 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 374642 0 374698 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 377770 0 377826 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 380806 0 380862 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 383842 0 383898 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 386878 0 386934 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 389914 0 389970 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 392950 0 393006 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 395986 0 396042 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 399022 0 399078 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 402058 0 402114 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 405094 0 405150 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 408130 0 408186 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 497808 6 vccd1
port 502 nsew power bidirectional
rlabel metal2 s 497738 499200 497794 500000 6 vccd1
port 503 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 497808 6 vssd1
port 504 nsew ground bidirectional
rlabel metal3 s 499200 249976 500000 250096 6 vssd1
port 505 nsew ground bidirectional
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 506 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 507 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 508 nsew signal output
rlabel metal2 s 6550 0 6606 800 6 wbs_adr_i[0]
port 509 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_adr_i[10]
port 510 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_adr_i[11]
port 511 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[12]
port 512 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[13]
port 513 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[14]
port 514 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[15]
port 515 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[16]
port 516 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 wbs_adr_i[17]
port 517 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_adr_i[18]
port 518 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_adr_i[19]
port 519 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[1]
port 520 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 wbs_adr_i[20]
port 521 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 wbs_adr_i[21]
port 522 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_adr_i[22]
port 523 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wbs_adr_i[23]
port 524 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[24]
port 525 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[25]
port 526 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 wbs_adr_i[26]
port 527 nsew signal input
rlabel metal2 s 92754 0 92810 800 6 wbs_adr_i[27]
port 528 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 wbs_adr_i[28]
port 529 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 wbs_adr_i[29]
port 530 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[2]
port 531 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 wbs_adr_i[30]
port 532 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_adr_i[31]
port 533 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[3]
port 534 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[4]
port 535 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_adr_i[5]
port 536 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[6]
port 537 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[7]
port 538 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_adr_i[8]
port 539 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[9]
port 540 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_cyc_i
port 541 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_dat_i[0]
port 542 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_dat_i[10]
port 543 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[11]
port 544 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_i[12]
port 545 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[13]
port 546 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_i[14]
port 547 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[15]
port 548 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[16]
port 549 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_dat_i[17]
port 550 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[18]
port 551 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_dat_i[19]
port 552 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_dat_i[1]
port 553 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wbs_dat_i[20]
port 554 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_i[21]
port 555 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_dat_i[22]
port 556 nsew signal input
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_i[23]
port 557 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[24]
port 558 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 wbs_dat_i[25]
port 559 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_i[26]
port 560 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_dat_i[27]
port 561 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_dat_i[28]
port 562 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[29]
port 563 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[2]
port 564 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 wbs_dat_i[30]
port 565 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wbs_dat_i[31]
port 566 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_i[3]
port 567 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_dat_i[4]
port 568 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[5]
port 569 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_i[6]
port 570 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_dat_i[7]
port 571 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_dat_i[8]
port 572 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[9]
port 573 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_o[0]
port 574 nsew signal output
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_o[10]
port 575 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[11]
port 576 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[12]
port 577 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[13]
port 578 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[14]
port 579 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_o[15]
port 580 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 wbs_dat_o[16]
port 581 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_o[17]
port 582 nsew signal output
rlabel metal2 s 67362 0 67418 800 6 wbs_dat_o[18]
port 583 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_o[19]
port 584 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[1]
port 585 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_o[20]
port 586 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 wbs_dat_o[21]
port 587 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[22]
port 588 nsew signal output
rlabel metal2 s 82542 0 82598 800 6 wbs_dat_o[23]
port 589 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wbs_dat_o[24]
port 590 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 wbs_dat_o[25]
port 591 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 wbs_dat_o[26]
port 592 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_o[27]
port 593 nsew signal output
rlabel metal2 s 97814 0 97870 800 6 wbs_dat_o[28]
port 594 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_o[29]
port 595 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[2]
port 596 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 wbs_dat_o[30]
port 597 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 wbs_dat_o[31]
port 598 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[3]
port 599 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_o[4]
port 600 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[5]
port 601 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_o[6]
port 602 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[7]
port 603 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[8]
port 604 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[9]
port 605 nsew signal output
rlabel metal2 s 9586 0 9642 800 6 wbs_sel_i[0]
port 606 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_sel_i[1]
port 607 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_sel_i[2]
port 608 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_sel_i[3]
port 609 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_stb_i
port 610 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_we_i
port 611 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 500000 500000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 247182584
string GDS_START 1472744
<< end >>

